library ieee;
use ieee.std_logic_1164.all;

entity writeback is

end writeback;

architecture rtl of writeback is

begin

end rtl;