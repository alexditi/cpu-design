library ieee;
use ieee.std_logic_1164.all;

library cpu_design;

entity cpu is

end cpu;

architecture rtl of cpu is

begin

end rtl;