library ieee;
use ieee.std_logic_1164.all;

library cpu_design;

entity cpu_embedded is

end cpu_embedded;

architecture rtl of cpu_embedded is

begin

end rtl;