library ieee;
use ieee.std_logic_1164.all;

entity and_gate is
	port (
		input_1    : in std_logic;
		input_2    : in std_logic;
		and_output : out std_logic
		);
end and_gate;

architecture rtl of and_gate is
	signal and_gate : std_logic;
begin
	and_gate <= input_1 and input_2;
	and_output <= and_gate;
end rtl;
